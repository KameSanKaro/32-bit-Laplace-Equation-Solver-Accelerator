--==============================================================================
--== Logisim-evolution goes FPGA automatic generated VHDL code                ==
--== https://github.com/logisim-evolution/                                    ==
--==                                                                          ==
--==                                                                          ==
--== Project   : Laplace32BitAccelerator-FPGA-TESTING                         ==
--== Component : synthesizedClockGenerator                                    ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY synthesizedClockGenerator IS
   PORT ( FPGAClock        : IN  std_logic;
          SynthesizedClock : OUT std_logic );
END ENTITY synthesizedClockGenerator;
